`timescale 1ns/1ps
`include "ALU.v"

module alu_test;

reg[31:0] instSet,reg_a,reg_b;
wire signed [31:0] res;
wire [2:0] flag;

alu test_alu(instSet, reg_a, reg_b, flag, res);

initial begin

    $dumpfile("output.vcd");
    $dumpvars(0, alu_test);

    $display("instruction:op:func:  reg_a   :  reg_b   :   RS   :  RT  : result : flag");
    $monitor("   %h:%h: %h :%h:%h:%h:%h:%h:%h",
    instSet, test_alu.opcode, test_alu.func, reg_a, reg_b, test_alu.RS, test_alu.RT, res, flag);

    // 1. add
    #10 instSet<=32'b0000_0000_0000_0000_0000_0000_0010_0000;
    reg_a<=32'b1000_0000_0000_0000_0000_0000_0000_0000;
    reg_b<=32'b1000_0000_0000_0000_0000_0000_0000_0000; 

    /*
    // 2. addi
    #10 instSet<=32'b0010_0000_0000_0000_0000_0000_0000_0001;
    reg_a <=32'b0000_0000_0000_0000_0000_0000_0000_0010;
    reg_b <= 32'b1000_0000_0000_0010_0000_0000_0001_0001;

    // 3. addu
    #10 instSet<=32'b0000_0000_0000_0000_0000_0000_0010_0001;
    reg_a<=32'b0000_0000_0000_0000_0000_0000_0000_0001;
    reg_b<=32'b0000_0000_0000_0000_0000_0000_0000_0010;

    // 4. addiu
    #10 instSet<=32'b0010_0100_0000_0000_0000_0000_0000_0001;
    reg_a<=32'b0000_0000_0000_0000_0000_0000_0000_0001;

    // 5. sub
    #10 instSet<=32'b0000_0000_0000_0000_0000_0000_0010_0010;
    reg_a<=32'b0000_0000_0000_0000_0000_0000_0000_0010;
    reg_b<=32'b0000_0000_0000_0000_0000_0000_0000_1010;

    // 6. subu
    #10 instSet<=32'b0000_0000_0000_0000_0000_0000_0010_0011;
    reg_a<=32'b0000_0000_0000_0000_0000_0000_0000_0010;
    reg_b<=32'b0000_0000_0000_0000_0000_0000_0000_0001;

    // 7. and
    #10 instSet<=32'b0000_0000_0000_0000_0000_0000_0010_0100;
    reg_a<=32'b0000_0000_0000_0000_0000_0000_0000_1001;
    reg_b<=32'b0000_0000_0000_0000_0000_0000_0000_1101;

    // 8. andi
    #10 instSet<=32'b0011_0000_0000_0000_0000_0000_0000_0001;
    reg_a<=32'b0000_0000_0000_0000_0000_0000_0000_1001;
    reg_b<= 32'b0000_0000_0000_0000_0000_0000_0000_0000;

    // 9. nor
    #10 instSet<=32'b0000_0000_0000_0000_0000_0000_0010_0111;
    reg_a<=32'b0000_0000_0000_0000_0000_0000_0000_1001;
    reg_b<=32'b0000_0000_0000_0000_0000_0000_0000_1101;

    // 10. or
    #10 instSet<=32'b0000_0000_0000_0000_0000_0000_0010_0101;
    reg_a<=32'b0000_0000_0000_0000_0000_0000_1001_0000;
    reg_b<=32'b0000_0000_0000_0000_0000_0000_1101_0000;

    // 11. ori
    #10 instSet<=32'b0011_0100_0000_0000_0000_0000_0000_1101;
    reg_a<=32'b0000_0000_0000_0000_0000_0000_0000_1001;
    reg_b<=32'b0000_0000_0000_0000_0000_0000_0000_0000;

    // 11. xor
    #10 instSet<=32'b0000_0000_0000_0000_0000_0000_0010_0110;
    reg_a<=32'b0000_0000_0000_0000_0000_0000_0000_1001;
    reg_b<=32'b0000_0000_0000_0000_0000_0000_0000_1101;

    // 13. xori
    #10 instSet<=32'b0011_1000_0000_0000_0000_0000_0000_1101;
    reg_a<=32'b0000_0000_0000_0000_0000_0000_0000_1001;
    reg_b<=32'b0000_0000_0000_0000_0000_0000_0000_0000;

    // 14. beq
    #10 instSet<=32'b0001_0000_0000_0000_0000_0000_0000_1000;
    reg_a<=32'b0000_0000_0000_0000_0000_0000_0000_1001;
    reg_b<=32'b0000_0000_0000_0000_0000_0000_0000_1001;

    // 15. bne
    #10 instSet<=32'b0001_0100_0000_0000_0000_0000_0000_1000;
    reg_a<=32'b0000_0000_0000_0000_0000_0000_0000_1001;
    reg_b<=32'b0000_0000_0000_0000_0000_0000_0000_1001;

    // 16. slt
    #10 instSet<=32'b0000_0000_0000_0001_0001_0000_0010_1010;
    reg_a<=32'b0000_0000_0000_0000_0000_0000_0000_1000;
    reg_b<=32'b0000_0000_0000_0000_0000_0000_0000_0001;

    // 17. slti
    #10 instSet<=32'b0010_1000_0000_0000_0000_0000_0000_1000;
    reg_a<=32'b0000_0000_0000_0000_0000_0000_0000_0001;

    // 18. sltiu
    #10 instSet<=32'b0010_1100_0000_0000_0000_0000_0000_1000;
    reg_a<=32'b0000_0000_0000_0000_0000_0000_0000_0001;

    // 19. sltu
    #10 instSet<=32'b0000_0000_0000_0000_0000_0000_0010_1011;
    reg_a<=32'b0000_0000_0000_0000_0000_0000_0000_0001;
    reg_b<=32'b0000_0000_0000_0000_0000_0000_0000_1000;

    // 20. lw
    #10 instSet<=32'b1000_1100_0000_0000_0000_0000_0000_1000;
    reg_b<=32'b0000_0000_0000_0000_0000_0000_0000_0000;

    // 21. sw
    #10 instSet<=32'b1010_1100_0000_0000_0000_0000_0000_0000;
    reg_a<=32'b0000_0000_0000_0000_0000_0000_0000_0000;
    reg_b<=32'b0000_0000_0000_0000_0000_0000_0000_1000;

    // 26. sll
    #10 instSet<=32'b0000_0000_0000_0000_0000_0000_0100_0000;
    reg_a<=32'b0000_0000_0000_0000_0000_0000_0000_0000;
    reg_b<=32'b1101_1101_1101_1101_1101_1101_1101_1101;

    // 27. sllv
    #10 instSet<=32'b0000_0000_0000_0000_0000_0000_0000_0100;
    reg_b<=32'b1101_1101_1101_1101_1101_1101_1101_1101;
    reg_a<=32'b0000_0000_0000_0000_0000_0000_0000_0100;

    // 28. srl
    #10 instSet<=32'b0000_0000_0000_0000_0000_0000_0000_0010;
    reg_a<=32'b0000_0000_0000_0000_0000_0000_0000_0100;
    reg_b<=32'b1101_1101_1101_1101_1101_1101_1101_1101;

    // 29. srlv
    #10 instSet<=32'b0000_0000_0000_0000_0000_0000_0000_0110;
    reg_b<=32'b1101_1101_1101_1101_1101_1101_1101_1101;
    reg_a<=32'b0000_0000_0000_0000_0000_0000_0000_0100;

    // 30. sra
    #10 instSet<=32'b0000_0000_0000_0000_0000_0000_0000_0011;
    reg_a <=32'b1101_1101_1101_1101_1101_1101_1101_1101;
    reg_b <=32'b0000_0000_0000_0000_0000_0000_0000_0000;

    // 31. srav
    #10 instSet<=32'b0000_0000_0000_0000_0000_0000_0000_0111;
    reg_b<=32'b1101_1101_1101_1101_1101_1101_1101_1101;
    reg_a<=32'b0000_0000_0000_0000_0000_0000_0000_0100;
    */

    #10 $finish;
    end
endmodule